`ifndef     INST_DEF
`define     INST_DEF

// 基础指令集青春版的机器码, 仅覆盖 alu, mdu, ls, branch 指令, 供 decoder 使用
`define     ADD     32'b0000_0000_0001_0000_0???_????_????_????
`define     SUB     32'b0000_0000_0001_0001_0???_????_????_????
`define     SLT     32'b0000_0000_0001_0010_0???_????_????_????
`define     SLTU    32'b0000_0000_0001_0010_1???_????_????_????
`define     NOR     32'b0000_0000_0001_0100_0???_????_????_????
`define     AND     32'b0000_0000_0001_0100_1???_????_????_????
`define     OR      32'b0000_0000_0001_0101_0???_????_????_????
`define     XOR     32'b0000_0000_0001_0101_1???_????_????_????
`define     SLL     32'b0000_0000_0001_0111_0???_????_????_????
`define     SRL     32'b0000_0000_0001_0111_1???_????_????_????
`define     SRA     32'b0000_0000_0001_1000_0???_????_????_????

`define     MUL     32'b0000_0000_0001_1100_0???_????_????_????
`define     MULH    32'b0000_0000_0001_1100_1???_????_????_????
`define     MULHU   32'b0000_0000_0001_1101_0???_????_????_????
`define     DIV     32'b0000_0000_0010_0000_0???_????_????_????
`define     MOD     32'b0000_0000_0010_0000_1???_????_????_????
`define     DIVU    32'b0000_0000_0010_0001_0???_????_????_????
`define     MODU    32'b0000_0000_0010_0001_1???_????_????_????

`define     SLLI    32'b0000_0000_0100_0000_1???_????_????_????
`define     SRLI    32'b0000_0000_0100_0100_1???_????_????_????
`define     SRAI    32'b0000_0000_0100_1000_1???_????_????_????

`define     SLTI    32'b0000_0010_00??_????_????_????_????_????
`define     SLTUI   32'b0000_0010_01??_????_????_????_????_????
`define     ADDI    32'b0000_0010_10??_????_????_????_????_????
`define     ANDI    32'b0000_0011_01??_????_????_????_????_????
`define     ORI     32'b0000_0011_10??_????_????_????_????_????
`define     SLTI    32'b0000_0011_11??_????_????_????_????_????

`define     LU12I   32'b0001_010?_????_????_????_????_????_????
`define     PCADD   32'b0001_110?_????_????_????_????_????_????

`define     LDB     32'b0010_1000_00??_????_????_????_????_????
`define     LDH     32'b0010_1000_01??_????_????_????_????_????
`define     LDW     32'b0010_1000_10??_????_????_????_????_????
`define     STB     32'b0010_1001_00??_????_????_????_????_????
`define     STH     32'b0010_1001_01??_????_????_????_????_????
`define     STW     32'b0010_1001_10??_????_????_????_????_????
`define     LDBU    32'b0010_1010_00??_????_????_????_????_????
`define     LDHU    32'b0010_1010_01??_????_????_????_????_????

// `define     JIRL    32'b0100_11??_????_????_????_????_????_????
`define     B       32'b0101_00??_????_????_????_????_????_????
`define     BL      32'b0101_01??_????_????_????_????_????_????
`define     BEQ     32'b0101_10??_????_????_????_????_????_????
`define     BNE     32'b0101_11??_????_????_????_????_????_????
`define     BLT     32'b0110_00??_????_????_????_????_????_????
`define     BGE     32'b0110_01??_????_????_????_????_????_????
`define     BLTU    32'b0110_10??_????_????_????_????_????_????
`define     BGEU    32'b0110_11??_????_????_????_????_????_????

`endif
