module PRF (
    input               clk,
    input               rst,
    input               stop,
    input               freeze_front,
    input               freeze_back,
    input               valid_issue,
    output              full_PRF,
    output  reg [4 : 0] tag_PRF,

    input       [4 : 0] tag_Ra_add,
    input       [4 : 0] tag_Rb_add,
    input       [4 : 0] tag_Ra_mul,
    input       [4 : 0] tag_Rb_mul,

    output      [15 : 0]busA_add,
    output      [15 : 0]busB_add,
    output      [15 : 0]busA_mul,
    output      [15 : 0]busB_mul,

    input               valid_Result_add,
    input       [15 : 0]Result_add,
    input       [4 : 0] tag_PRF_add,
    input               valid_Result_mul,
    input       [15 : 0]Result_mul,
    input       [4 : 0] tag_PRF_mul,

    input       [4 : 0] ARF_tag [7 : 0],
    input               RegWr_ARF,
    input       [4 : 0] tag_PRF_ARF,
    input       [4 : 0] tag_Rw_old
);

    reg     [15 : 0]    data [31 : 0];
    reg     [31 : 0]    free_list;

    integer i;

    always @(posedge clk or negedge rst) begin
        if (!rst) begin
            for (i = 0; i < 32; i = i + 1) begin
                data[i] <= i;
            end
            free_list <= 32'hffff_ff00;
        end
        else if (!stop) begin
            if (!freeze_front && valid_issue) begin
                free_list[tag_PRF] <= 0;
            end
            if (!freeze_back && valid_Result_add && tag_PRF_add != 0) begin
                data[tag_PRF_add] <= Result_add;
            end
            if (!freeze_back && valid_Result_mul && tag_PRF_mul != 0) begin
                data[tag_PRF_mul] <= Result_mul;
            end
            if (RegWr_ARF && tag_PRF_ARF != 0) begin
                free_list[tag_Rw_old] <= 1;
            end
        end
        else begin
            free_list <= 32'hffff_ffff;
            for (i = 0; i < 8; i = i + 1) begin
                free_list[ARF_tag[i]] <= 0;
            end
        end
    end

    always @(*) begin
        casez (free_list)
            32'b????_????_????_????_????_????_????_???1:    tag_PRF = 0;
            32'b????_????_????_????_????_????_????_??10:    tag_PRF = 1;
            32'b????_????_????_????_????_????_????_?100:    tag_PRF = 2;
            32'b????_????_????_????_????_????_????_1000:    tag_PRF = 3;
            32'b????_????_????_????_????_????_???1_0000:    tag_PRF = 4;
            32'b????_????_????_????_????_????_??10_0000:    tag_PRF = 5;
            32'b????_????_????_????_????_????_?100_0000:    tag_PRF = 6;
            32'b????_????_????_????_????_????_1000_0000:    tag_PRF = 7;

            32'b????_????_????_????_????_???1_0000_0000:    tag_PRF = 8;
            32'b????_????_????_????_????_??10_0000_0000:    tag_PRF = 9;
            32'b????_????_????_????_????_?100_0000_0000:    tag_PRF = 10;
            32'b????_????_????_????_????_1000_0000_0000:    tag_PRF = 11;
            32'b????_????_????_????_???1_0000_0000_0000:    tag_PRF = 12;
            32'b????_????_????_????_??10_0000_0000_0000:    tag_PRF = 13;
            32'b????_????_????_????_?100_0000_0000_0000:    tag_PRF = 14;
            32'b????_????_????_????_1000_0000_0000_0000:    tag_PRF = 15;

            32'b????_????_????_???1_0000_0000_0000_0000:    tag_PRF = 16;
            32'b????_????_????_??10_0000_0000_0000_0000:    tag_PRF = 17;
            32'b????_????_????_?100_0000_0000_0000_0000:    tag_PRF = 18;
            32'b????_????_????_1000_0000_0000_0000_0000:    tag_PRF = 19;
            32'b????_????_???1_0000_0000_0000_0000_0000:    tag_PRF = 20;
            32'b????_????_??10_0000_0000_0000_0000_0000:    tag_PRF = 21;
            32'b????_????_?100_0000_0000_0000_0000_0000:    tag_PRF = 22;
            32'b????_????_1000_0000_0000_0000_0000_0000:    tag_PRF = 23;

            32'b????_???1_0000_0000_0000_0000_0000_0000:    tag_PRF = 24;
            32'b????_??10_0000_0000_0000_0000_0000_0000:    tag_PRF = 25;
            32'b????_?100_0000_0000_0000_0000_0000_0000:    tag_PRF = 26;
            32'b????_1000_0000_0000_0000_0000_0000_0000:    tag_PRF = 27;
            32'b???1_0000_0000_0000_0000_0000_0000_0000:    tag_PRF = 28;
            32'b??10_0000_0000_0000_0000_0000_0000_0000:    tag_PRF = 29;
            32'b?100_0000_0000_0000_0000_0000_0000_0000:    tag_PRF = 30;
            32'b1000_0000_0000_0000_0000_0000_0000_0000:    tag_PRF = 31;
            default:                                        tag_PRF = 0;
        endcase
    end

    assign  full_PRF = (free_list == 32'h0000_0000)? 1 : 0;
    
    assign  busA_add = data[tag_Ra_add];
    assign  busB_add = data[tag_Rb_add];
    assign  busA_mul = data[tag_Ra_mul];
    assign  busB_mul = data[tag_Rb_mul];

endmodule