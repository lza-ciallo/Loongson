module IM (
    input clk,
    input rst,
    input [31:0] pc,
    output [31:0] inst[2:0],
    output inst_valid[2:0]
);
endmodule
