module IF_ID (
    // IF SIGNALS


    // ID SIGNALS


    // s
);

endmodule
