module SRAT (
    input               clk,
    input               rst,
    input               freeze_front,
    input               valid_pc,
    output              full_PRF,
    // x,y,z 端口读写
    input   [ 1 : 0]    Type        [2 : 0],
    input   [ 2 : 0]    Ra          [2 : 0],
    input   [ 2 : 0]    Rb          [2 : 0],
    input   [ 2 : 0]    Rw          [2 : 0],
    output  [ 4 : 0]    Pa          [2 : 0],
    output  [ 4 : 0]    Pb          [2 : 0],
    output  [ 4 : 0]    Pw          [2 : 0],
    output  [ 4 : 0]    Pw_old      [2 : 0],
    output              valid_Pa    [2 : 0],
    output              valid_Pb    [2 : 0],
    // ADD 广播
    input   [ 4 : 0]    Pw_Result_add,
    input               valid_Result_add,
    // MUL 广播
    input   [ 4 : 0]    Pw_Result_mul,
    input               valid_Result_mul,
    // LS 广播
    input   [ 4 : 0]    Pw_Result_ls,
    input               valid_Result_ls,
    input               mode_ls,    // 1 为写, 0 为读
    // ROB 退休
    input               ready_ret   [2 : 0],
    input               excep_ret   [2 : 0],
    input   [ 1 : 0]    Type_ret    [2 : 0],
    input   [ 4 : 0]    Pw_old_ret  [2 : 0],
    // 精确异常恢复
    input               flush,
    input   [ 4 : 0]    ARAT_P_list [7 : 0],
    input   [31 : 0]    ARAT_freelist
);

    // typedef struct packed {
    //     reg [ 4 : 0]    P_list;
    //     reg             valid_list;
    // } srat_list;

    // srat_list           list    [7 : 0];

    reg     [ 4 : 0]    P_list  [7 : 0];    // +
    reg     [31 : 0]    valid_list;         // +

    reg     [ 4 : 0]    Pw_r    [2 : 0];

    reg     [31 : 0]    free_list;
    wire    [31 : 0]    free_list_y;
    wire    [31 : 0]    free_list_z;

    integer i;

    // 写入 Pw, 接收广播, ROB 退休释放
    always @(posedge clk or negedge rst) begin
        if (!rst) begin
            for (i = 0; i < 8; i = i + 1) begin
                // list[i].P_list      <=  i;
                // list[i].valid_list  <=  1;
                P_list[i]   <=  i;          // +
            end
            valid_list  <=  32'h0000_00ff;  // +
            free_list   <=  32'hffff_ff00;
        end
        else begin
            if (!flush) begin
                
                // 前端记录新分配的 Rw-Pw
                if (valid_pc && !freeze_front) begin
                    if (Type[0] != 2'b11) begin
                        free_list[Pw[0]]    <=  0;
                        if (Rw[0] != 0 && !((Type[1] != 2'b11 && Rw[0] == Rw[1]) || (Type[2] != 2'b11 && Rw[0] == Rw[2]))) begin
                            // list[Rw[0]]     <=  {Pw[0], 1'b0};
                            P_list[Rw[0]]       <=  Pw[0];  // +
                            valid_list[Pw[0]]   <=  0;      // +
                        end
                    end
                    if (Type[1] != 2'b11) begin
                        free_list[Pw[1]]    <=  0;
                        if (Rw[1] != 0 && !(Type[2] != 2'b11 && Rw[1] == Rw[2])) begin
                            // list[Rw[1]]     <=  {Pw[1], 1'b0};
                            P_list[Rw[1]]       <=  Pw[1];  // +
                            valid_list[Pw[1]]   <=  0;      // +
                        end
                    end
                    if (Type[2] != 2'b11) begin
                        free_list[Pw[2]]    <=  0;
                        if (Rw[2] != 0) begin
                            // list[Rw[2]]     <=  {Pw[2], 1'b0};
                            P_list[Rw[2]]       <=  Pw[2];  // +
                            valid_list[Pw[2]]   <=  0;      // +
                        end
                    end
                end

                // 接收广播信号
                if (valid_Result_add) begin
                    // for (i = 0; i < 8; i = i + 1) begin
                    //     if (!(valid_pc && !freeze_front &&
                    //         ((i == Rw[0] && Type[0] != 2'b11) || (i == Rw[1] && Type[1] != 2'b11) || (i == Rw[1] && Type[1] != 2'b11)))) begin
                    //         if (list[i].P_list == Pw_Result_add) begin
                    //             list[i].valid_list <= 1;
                    //         end
                    //     end
                    // end
                    valid_list[Pw_Result_add]   <=  1;  // +
                end
                if (valid_Result_mul) begin
                    // for (i = 0; i < 8; i = i + 1) begin
                    //     if (!(valid_pc && !freeze_front &&
                    //         ((i == Rw[0] && Type[0] != 2'b11) || (i == Rw[1] && Type[1] != 2'b11) || (i == Rw[1] && Type[1] != 2'b11)))) begin
                    //         if (list[i].P_list == Pw_Result_mul) begin
                    //             list[i].valid_list <= 1;
                    //         end
                    //     end
                    // end
                    valid_list[Pw_Result_mul]   <=  1;  // +
                end
                if (valid_Result_ls && mode_ls == 1) begin
                    // for (i = 0; i < 8; i = i + 1) begin
                    //     if (!(valid_pc && !freeze_front &&
                    //         ((i == Rw[0] && Type[0] != 2'b11) || (i == Rw[1] && Type[1] != 2'b11) || (i == Rw[1] && Type[1] != 2'b11)))) begin
                    //         if (list[i].P_list == Pw_Result_ls) begin
                    //             list[i].valid_list <= 1;
                    //         end
                    //     end
                    // end
                    valid_list[Pw_Result_ls]    <=  1;  // +
                end

                // 退休后释放 free_list
                if (ready_ret[0] && !excep_ret[0]) begin
                    if (Pw_old_ret[0] != 0) begin
                        free_list[Pw_old_ret[0]] <= 1;
                    end
                    if (ready_ret[1] && !excep_ret[1]) begin
                        if (Pw_old_ret[1] != 0) begin
                            free_list[Pw_old_ret[1]] <= 1;
                        end
                        if (ready_ret[2] && !excep_ret[2]) begin
                            if (Pw_old_ret[2] != 0) begin
                                free_list[Pw_old_ret[2]] <= 1;
                            end
                        end
                    end
                end
            end

            // 精确异常恢复
            else begin
                // for (i = 0; i < 8; i = i + 1) begin
                    // list[i] <=  {ARAT_P_list[i], 1'b1};
                // end
                P_list      <=  ARAT_P_list;        // +
                valid_list  <=  ~ARAT_freelist;     // +
                free_list   <=  ARAT_freelist;
            end
        end
    end

    // x,y,z 端口读 Pa,Pb,Pw_old
    // assign  {Pa[0], valid_Pa[0]}    =   list[Ra[0]];
    // assign  {Pb[0], valid_Pb[0]}    =   list[Rb[0]];
    // assign  Pw_old[0]               =   list[Rw[0]].P_list;

    // assign  {Pa[1], valid_Pa[1]}    =   (Ra[1] == 0)? list[Ra[1]] : (Ra[1] == Rw[0])? {Pw[0], 1'b0} : list[Ra[1]];
    // assign  {Pb[1], valid_Pb[1]}    =   (Rb[1] == 0)? list[Rb[1]] : (Rb[1] == Rw[0])? {Pw[0], 1'b0} : list[Rb[1]];
    // assign  Pw_old[1]               =                               (Rw[1] == Rw[0])? Pw[0]         : list[Rw[1]].P_list;

    // assign  {Pa[2], valid_Pa[2]}    =   (Ra[2] == 0)? list[Ra[2]] : (Ra[2] == Rw[1])? {Pw[1], 1'b0} :
    //                                                                 (Ra[2] == Rw[0])? {Pw[0], 1'b0} : list[Ra[2]];
    // assign  {Pb[2], valid_Pb[2]}    =   (Rb[2] == 0)? list[Rb[2]] : (Rb[2] == Rw[1])? {Pw[1], 1'b0} :
    //                                                                 (Rb[2] == Rw[0])? {Pw[0], 1'b0} : list[Rb[2]];
    // assign  Pw_old[2]               =                               (Rw[2] == Rw[1])? Pw[1]         :
    //                                                                 (Rw[2] == Rw[0])? Pw[0]         : list[Rw[2]].P_list;

    // +
    assign  Pa[0]       =   P_list[Ra[0]];
    assign  Pb[0]       =   P_list[Rb[0]];
    assign  Pw_old[0]   =   P_list[Rw[0]];
    assign  valid_Pa[0] =   valid_list[Pa[0]];
    assign  valid_Pb[0] =   valid_list[Pb[0]];

    assign  Pa[1]       =   (Ra[1] == 0)? P_list[Ra[1]] :   (Ra[1] == Rw[0])? Pw[0] : P_list[Ra[1]];
    assign  Pb[1]       =   (Rb[1] == 0)? P_list[Rb[1]] :   (Rb[1] == Rw[0])? Pw[0] : P_list[Rb[1]];
    assign  Pw_old[1]   =                                   (Rw[1] == Rw[0])? Pw[0] : P_list[Rw[1]];
    assign  valid_Pa[1] =   (Ra[1] == 0)? 1             :   (Ra[1] == Rw[0])? 0     : valid_list[Pa[1]];
    assign  valid_Pb[1] =   (Rb[1] == 0)? 1             :   (Rb[1] == Rw[0])? 0     : valid_list[Pb[1]];

    assign  Pa[2]       =   (Ra[2] == 0)? P_list[Ra[2]] :   (Ra[2] == Rw[1])? Pw[1] :
                                                            (Ra[2] == Rw[0])? Pw[0] : P_list[Ra[2]];
    assign  Pb[2]       =   (Rb[2] == 0)? P_list[Rb[2]] :   (Rb[2] == Rw[1])? Pw[1] :
                                                            (Rb[2] == Rw[0])? Pw[0] : P_list[Rb[2]];
    assign  Pw_old[2]   =                                   (Rw[2] == Rw[1])? Pw[1] :
                                                            (Rw[2] == Rw[0])? Pw[0] : P_list[Rw[2]];
    assign  valid_Pa[2] =   (Ra[2] == 0)? 1             :   (Ra[2] == Rw[1])? 0     :
                                                            (Ra[2] == Rw[0])? 0     : valid_list[Pa[2]];
    assign  valid_Pb[2] =   (Rb[2] == 0)? 1             :   (Rb[2] == Rw[1])? 0     :
                                                            (Rb[2] == Rw[0])? 0     : valid_list[Pb[2]];
    // +

    // 分配 Pw, 并生成 full_PRF
    assign  Pw[0]   =   (Rw[0] == 0)? 0 : Pw_r[0];
    assign  Pw[1]   =   (Rw[1] == 0)? 0 : Pw_r[1];
    assign  Pw[2]   =   (Rw[2] == 0)? 0 : Pw_r[2];

    assign  free_list_y =   free_list   &   ~(32'd1 << Pw[0]);
    assign  free_list_z =   free_list_y &   ~(32'd1 << Pw[1]);

    assign  full_PRF_x  = (free_list    ==  32'd0)? 1 : 0;
    assign  full_PRF_y  = (free_list_y  ==  32'd0)? 1 : 0;
    assign  full_PRF_z  = (free_list_z  ==  32'd0)? 1 : 0;
    assign  full_PRF    = (full_PRF_x || full_PRF_y || full_PRF_z)? 1 : 0;

    always @(*) begin
        // 端口 x 分配 (Pw_r[0])
        casez (free_list)
            32'b????_????_????_????_????_????_????_???1:    Pw_r[0] = 5'd0;
            32'b????_????_????_????_????_????_????_??10:    Pw_r[0] = 5'd1;
            32'b????_????_????_????_????_????_????_?100:    Pw_r[0] = 5'd2;
            32'b????_????_????_????_????_????_????_1000:    Pw_r[0] = 5'd3;
            32'b????_????_????_????_????_????_???1_0000:    Pw_r[0] = 5'd4;
            32'b????_????_????_????_????_????_??10_0000:    Pw_r[0] = 5'd5;
            32'b????_????_????_????_????_????_?100_0000:    Pw_r[0] = 5'd6;
            32'b????_????_????_????_????_????_1000_0000:    Pw_r[0] = 5'd7;

            32'b????_????_????_????_????_???1_0000_0000:    Pw_r[0] = 5'd8;
            32'b????_????_????_????_????_??10_0000_0000:    Pw_r[0] = 5'd9;
            32'b????_????_????_????_????_?100_0000_0000:    Pw_r[0] = 5'd10;
            32'b????_????_????_????_????_1000_0000_0000:    Pw_r[0] = 5'd11;
            32'b????_????_????_????_???1_0000_0000_0000:    Pw_r[0] = 5'd12;
            32'b????_????_????_????_??10_0000_0000_0000:    Pw_r[0] = 5'd13;
            32'b????_????_????_????_?100_0000_0000_0000:    Pw_r[0] = 5'd14;
            32'b????_????_????_????_1000_0000_0000_0000:    Pw_r[0] = 5'd15;

            32'b????_????_????_???1_0000_0000_0000_0000:    Pw_r[0] = 5'd16;
            32'b????_????_????_??10_0000_0000_0000_0000:    Pw_r[0] = 5'd17;
            32'b????_????_????_?100_0000_0000_0000_0000:    Pw_r[0] = 5'd18;
            32'b????_????_????_1000_0000_0000_0000_0000:    Pw_r[0] = 5'd19;
            32'b????_????_???1_0000_0000_0000_0000_0000:    Pw_r[0] = 5'd20;
            32'b????_????_??10_0000_0000_0000_0000_0000:    Pw_r[0] = 5'd21;
            32'b????_????_?100_0000_0000_0000_0000_0000:    Pw_r[0] = 5'd22;
            32'b????_????_1000_0000_0000_0000_0000_0000:    Pw_r[0] = 5'd23;

            32'b????_???1_0000_0000_0000_0000_0000_0000:    Pw_r[0] = 5'd24;
            32'b????_??10_0000_0000_0000_0000_0000_0000:    Pw_r[0] = 5'd25;
            32'b????_?100_0000_0000_0000_0000_0000_0000:    Pw_r[0] = 5'd26;
            32'b????_1000_0000_0000_0000_0000_0000_0000:    Pw_r[0] = 5'd27;
            32'b???1_0000_0000_0000_0000_0000_0000_0000:    Pw_r[0] = 5'd28;
            32'b??10_0000_0000_0000_0000_0000_0000_0000:    Pw_r[0] = 5'd29;
            32'b?100_0000_0000_0000_0000_0000_0000_0000:    Pw_r[0] = 5'd30;
            32'b1000_0000_0000_0000_0000_0000_0000_0000:    Pw_r[0] = 5'd31;
            default:                                        Pw_r[0] = 5'd0;
        endcase

        // 端口 y 分配 (Pw_r[1])
        casez (free_list_y)
            32'b????_????_????_????_????_????_????_???1:    Pw_r[1] = 5'd0;
            32'b????_????_????_????_????_????_????_??10:    Pw_r[1] = 5'd1;
            32'b????_????_????_????_????_????_????_?100:    Pw_r[1] = 5'd2;
            32'b????_????_????_????_????_????_????_1000:    Pw_r[1] = 5'd3;
            32'b????_????_????_????_????_????_???1_0000:    Pw_r[1] = 5'd4;
            32'b????_????_????_????_????_????_??10_0000:    Pw_r[1] = 5'd5;
            32'b????_????_????_????_????_????_?100_0000:    Pw_r[1] = 5'd6;
            32'b????_????_????_????_????_????_1000_0000:    Pw_r[1] = 5'd7;

            32'b????_????_????_????_????_???1_0000_0000:    Pw_r[1] = 5'd8;
            32'b????_????_????_????_????_??10_0000_0000:    Pw_r[1] = 5'd9;
            32'b????_????_????_????_????_?100_0000_0000:    Pw_r[1] = 5'd10;
            32'b????_????_????_????_????_1000_0000_0000:    Pw_r[1] = 5'd11;
            32'b????_????_????_????_???1_0000_0000_0000:    Pw_r[1] = 5'd12;
            32'b????_????_????_????_??10_0000_0000_0000:    Pw_r[1] = 5'd13;
            32'b????_????_????_????_?100_0000_0000_0000:    Pw_r[1] = 5'd14;
            32'b????_????_????_????_1000_0000_0000_0000:    Pw_r[1] = 5'd15;

            32'b????_????_????_???1_0000_0000_0000_0000:    Pw_r[1] = 5'd16;
            32'b????_????_????_??10_0000_0000_0000_0000:    Pw_r[1] = 5'd17;
            32'b????_????_????_?100_0000_0000_0000_0000:    Pw_r[1] = 5'd18;
            32'b????_????_????_1000_0000_0000_0000_0000:    Pw_r[1] = 5'd19;
            32'b????_????_???1_0000_0000_0000_0000_0000:    Pw_r[1] = 5'd20;
            32'b????_????_??10_0000_0000_0000_0000_0000:    Pw_r[1] = 5'd21;
            32'b????_????_?100_0000_0000_0000_0000_0000:    Pw_r[1] = 5'd22;
            32'b????_????_1000_0000_0000_0000_0000_0000:    Pw_r[1] = 5'd23;

            32'b????_???1_0000_0000_0000_0000_0000_0000:    Pw_r[1] = 5'd24;
            32'b????_??10_0000_0000_0000_0000_0000_0000:    Pw_r[1] = 5'd25;
            32'b????_?100_0000_0000_0000_0000_0000_0000:    Pw_r[1] = 5'd26;
            32'b????_1000_0000_0000_0000_0000_0000_0000:    Pw_r[1] = 5'd27;
            32'b???1_0000_0000_0000_0000_0000_0000_0000:    Pw_r[1] = 5'd28;
            32'b??10_0000_0000_0000_0000_0000_0000_0000:    Pw_r[1] = 5'd29;
            32'b?100_0000_0000_0000_0000_0000_0000_0000:    Pw_r[1] = 5'd30;
            32'b1000_0000_0000_0000_0000_0000_0000_0000:    Pw_r[1] = 5'd31;
            default:                                        Pw_r[1] = 5'd0;
        endcase

        // 端口 z 分配 (Pw_r[2])
        casez (free_list_z)
            32'b????_????_????_????_????_????_????_???1:    Pw_r[2] = 5'd0;
            32'b????_????_????_????_????_????_????_??10:    Pw_r[2] = 5'd1;
            32'b????_????_????_????_????_????_????_?100:    Pw_r[2] = 5'd2;
            32'b????_????_????_????_????_????_????_1000:    Pw_r[2] = 5'd3;
            32'b????_????_????_????_????_????_???1_0000:    Pw_r[2] = 5'd4;
            32'b????_????_????_????_????_????_??10_0000:    Pw_r[2] = 5'd5;
            32'b????_????_????_????_????_????_?100_0000:    Pw_r[2] = 5'd6;
            32'b????_????_????_????_????_????_1000_0000:    Pw_r[2] = 5'd7;

            32'b????_????_????_????_????_???1_0000_0000:    Pw_r[2] = 5'd8;
            32'b????_????_????_????_????_??10_0000_0000:    Pw_r[2] = 5'd9;
            32'b????_????_????_????_????_?100_0000_0000:    Pw_r[2] = 5'd10;
            32'b????_????_????_????_????_1000_0000_0000:    Pw_r[2] = 5'd11;
            32'b????_????_????_????_???1_0000_0000_0000:    Pw_r[2] = 5'd12;
            32'b????_????_????_????_??10_0000_0000_0000:    Pw_r[2] = 5'd13;
            32'b????_????_????_????_?100_0000_0000_0000:    Pw_r[2] = 5'd14;
            32'b????_????_????_????_1000_0000_0000_0000:    Pw_r[2] = 5'd15;

            32'b????_????_????_???1_0000_0000_0000_0000:    Pw_r[2] = 5'd16;
            32'b????_????_????_??10_0000_0000_0000_0000:    Pw_r[2] = 5'd17;
            32'b????_????_????_?100_0000_0000_0000_0000:    Pw_r[2] = 5'd18;
            32'b????_????_????_1000_0000_0000_0000_0000:    Pw_r[2] = 5'd19;
            32'b????_????_???1_0000_0000_0000_0000_0000:    Pw_r[2] = 5'd20;
            32'b????_????_??10_0000_0000_0000_0000_0000:    Pw_r[2] = 5'd21;
            32'b????_????_?100_0000_0000_0000_0000_0000:    Pw_r[2] = 5'd22;
            32'b????_????_1000_0000_0000_0000_0000_0000:    Pw_r[2] = 5'd23;

            32'b????_???1_0000_0000_0000_0000_0000_0000:    Pw_r[2] = 5'd24;
            32'b????_??10_0000_0000_0000_0000_0000_0000:    Pw_r[2] = 5'd25;
            32'b????_?100_0000_0000_0000_0000_0000_0000:    Pw_r[2] = 5'd26;
            32'b????_1000_0000_0000_0000_0000_0000_0000:    Pw_r[2] = 5'd27;
            32'b???1_0000_0000_0000_0000_0000_0000_0000:    Pw_r[2] = 5'd28;
            32'b??10_0000_0000_0000_0000_0000_0000_0000:    Pw_r[2] = 5'd29;
            32'b?100_0000_0000_0000_0000_0000_0000_0000:    Pw_r[2] = 5'd30;
            32'b1000_0000_0000_0000_0000_0000_0000_0000:    Pw_r[2] = 5'd31;
            default:                                        Pw_r[2] = 5'd0;
        endcase
    end

endmodule