module SRAT (
    input               clk,
    input               rst,
    input               freeze_front,
    output              full_PRF,
    // 端口 x 读写
    input               valid_issue_x,
    input   [2 : 0]     Ra_x,
    input   [2 : 0]     Rb_x,
    input   [2 : 0]     Rw_x,
    output  [4 : 0]     Pw_x,
    output  [4 : 0]     Pa_x,
    output  [4 : 0]     Pb_x,
    output  [4 : 0]     Pw_old_x,
    output              valid_Ra_x,
    output              valid_Rb_x,
    // 端口 y 读写
    input               valid_issue_y,
    input   [2 : 0]     Ra_y,
    input   [2 : 0]     Rb_y,
    input   [2 : 0]     Rw_y,
    output  [4 : 0]     Pw_y,
    output  [4 : 0]     Pa_y,
    output  [4 : 0]     Pb_y,
    output  [4 : 0]     Pw_old_y,
    output              valid_Ra_y,
    output              valid_Rb_y,
    // 端口 z 读写
    input               valid_issue_z,
    input   [2 : 0]     Ra_z,
    input   [2 : 0]     Rb_z,
    input   [2 : 0]     Rw_z,
    output  [4 : 0]     Pw_z,
    output  [4 : 0]     Pa_z,
    output  [4 : 0]     Pb_z,
    output  [4 : 0]     Pw_old_z,
    output              valid_Ra_z,
    output              valid_Rb_z,
    // 广播
    input   [4 : 0]     Pw_Result_add,
    input               valid_Result_add,
    input   [4 : 0]     Pw_Result_mul,
    input               valid_Result_mul,
    // ROB 退休释放 free_list
    input               RegWr_x,
    input               RegWr_y,
    input               RegWr_z,
    input               exp_x,
    input               exp_y,
    input               exp_z,
    input   [4 : 0]     Pw_retire_x,
    input   [4 : 0]     Pw_retire_y,
    input   [4 : 0]     Pw_retire_z,
    // 精确异常恢复
    input               flush,
    input   [4 : 0]     ARAT_P_list [7 : 0]
);

    reg     [4 : 0]     Pw_x_r;
    reg     [4 : 0]     Pw_y_r;
    reg     [4 : 0]     Pw_z_r;
    
    assign  Pw_x = (Rw_x == 0)? 0 : Pw_x_r;
    assign  Pw_y = (Rw_y == 0)? 0 : Pw_y_r;
    assign  Pw_z = (Rw_z == 0)? 0 : Pw_z_r;

    reg     [7 : 0]     valid_list;
    reg     [31 : 0]    free_list;
    reg     [4 : 0]     P_list [7 : 0];

    wire    [31 : 0]    free_list_y;
    wire    [31 : 0]    free_list_z;

    assign  Pa_x = P_list[Ra_x];
    assign  Pb_x = P_list[Rb_x];
    assign  Pw_old_x = P_list[Rw_x];
    assign  valid_Ra_x = valid_list[Ra_x];
    assign  valid_Rb_x = valid_list[Rb_x];

    assign  Pa_y = (Ra_y == Rw_x)? Pw_x : P_list[Ra_y];
    assign  Pb_y = (Rb_y == Rw_x)? Pw_x : P_list[Rb_y];
    assign  Pw_old_y = (Rw_y == Rw_x)? Pw_x : P_list[Rw_y];
    assign  valid_Ra_y = (Ra_y == Rw_x)? 0 : valid_list[Ra_y];
    assign  valid_Rb_y = (Rb_y == Rw_x)? 0 : valid_list[Rb_y];

    assign  Pa_z = (Ra_z == Rw_y)? Pw_y : (Ra_z == Rw_x)? Pw_x : P_list[Ra_z];
    assign  Pb_z = (Rb_z == Rw_y)? Pw_y : (Rb_z == Rw_x)? Pw_x : P_list[Rb_z];
    assign  Pw_old_z = (Rw_z == Rw_y)? Pw_y : (Rw_z == Rw_x)? Pw_x : P_list[Rw_z];
    assign  valid_Ra_z = (Ra_z == Rw_y || Ra_z == Rw_x)? 0 : valid_list[Ra_z];
    assign  valid_Rb_z = (Rb_z == Rw_y || Rb_z == Rw_x)? 0 : valid_list[Rb_z];

    integer i;

    always @(posedge clk or negedge rst) begin
        if (!rst) begin
            valid_list <= 8'hff;
            free_list <= 32'hffff_ff00;
            for (i = 0; i < 8; i = i + 1) begin
                P_list[i] <= i;
            end
        end
        else begin
            if (!flush) begin
                // 前端记录新分配的 Rw-Pw
                if (!freeze_front) begin
                    if (valid_issue_x) begin
                        free_list[Pw_x] <= 0;
                        if (Rw_x != 0 && !((valid_issue_y && Rw_x == Rw_y) || (valid_issue_z && Rw_x == Rw_z))) begin
                            valid_list[Rw_x] <= 0;
                            P_list[Rw_x] <= Pw_x;
                        end
                    end
                    if (valid_issue_y) begin
                        free_list[Pw_y] <= 0;
                        if (Rw_y != 0 && !(valid_issue_z && Rw_y == Rw_z)) begin
                            valid_list[Rw_y] <= 0;
                            P_list[Rw_y] <= Pw_y;
                        end
                    end
                    if (valid_issue_z) begin
                        free_list[Pw_z] <= 0;
                        if (Rw_z != 0) begin
                            valid_list[Rw_z] <= 0;
                            P_list[Rw_z] <= Pw_z;
                        end
                    end
                end
                // 接收广播信号
                if (valid_Result_add) begin
                    for (i = 0; i < 8; i = i + 1) begin
                        if ((i != Rw_x && i != Rw_y && i != Rw_z) || freeze_front ||
                            (!valid_issue_x && !valid_issue_y && !valid_issue_z)) begin
                            if (P_list[i] == Pw_Result_add) begin
                                valid_list[i] <= 1;
                            end
                        end
                    end
                end
                if (valid_Result_mul) begin
                    for (i = 0; i < 8; i = i + 1) begin
                        if ((i != Rw_x && i != Rw_y && i != Rw_z) || freeze_front ||
                            (!valid_issue_x && !valid_issue_y && !valid_issue_z)) begin
                            if (P_list[i] == Pw_Result_mul) begin
                                valid_list[i] <= 1;
                            end
                        end
                    end
                end
                // 退休后释放 free_list
                if (RegWr_x && !exp_x) begin
                    free_list[Pw_retire_x] <= 1;
                    if (RegWr_y && !exp_y) begin
                        free_list[Pw_retire_y] <= 1;
                        if (RegWr_z && !exp_z) begin
                            free_list[Pw_retire_z] <= 1;
                        end
                    end
                end
            end
            // 精确异常恢复
            else begin
                P_list <= ARAT_P_list;
                valid_list <= 8'hff;
                free_list <= 32'hffff_ffff;
                for (i = 0; i < 8; i = i + 1) begin
                    free_list[ARAT_P_list[i]] <= 0;
                end
            end
        end
    end

    assign  free_list_y = free_list & ~(32'd1 << Pw_x);
    assign  free_list_z = free_list_y & ~(32'd1 << Pw_y);

    always @(*) begin
       casez (free_list)
            32'b????_????_????_????_????_????_????_???1:    Pw_x_r = 0;
            32'b????_????_????_????_????_????_????_??10:    Pw_x_r = 1;
            32'b????_????_????_????_????_????_????_?100:    Pw_x_r = 2;
            32'b????_????_????_????_????_????_????_1000:    Pw_x_r = 3;
            32'b????_????_????_????_????_????_???1_0000:    Pw_x_r = 4;
            32'b????_????_????_????_????_????_??10_0000:    Pw_x_r = 5;
            32'b????_????_????_????_????_????_?100_0000:    Pw_x_r = 6;
            32'b????_????_????_????_????_????_1000_0000:    Pw_x_r = 7;

            32'b????_????_????_????_????_???1_0000_0000:    Pw_x_r = 8;
            32'b????_????_????_????_????_??10_0000_0000:    Pw_x_r = 9;
            32'b????_????_????_????_????_?100_0000_0000:    Pw_x_r = 10;
            32'b????_????_????_????_????_1000_0000_0000:    Pw_x_r = 11;
            32'b????_????_????_????_???1_0000_0000_0000:    Pw_x_r = 12;
            32'b????_????_????_????_??10_0000_0000_0000:    Pw_x_r = 13;
            32'b????_????_????_????_?100_0000_0000_0000:    Pw_x_r = 14;
            32'b????_????_????_????_1000_0000_0000_0000:    Pw_x_r = 15;

            32'b????_????_????_???1_0000_0000_0000_0000:    Pw_x_r = 16;
            32'b????_????_????_??10_0000_0000_0000_0000:    Pw_x_r = 17;
            32'b????_????_????_?100_0000_0000_0000_0000:    Pw_x_r = 18;
            32'b????_????_????_1000_0000_0000_0000_0000:    Pw_x_r = 19;
            32'b????_????_???1_0000_0000_0000_0000_0000:    Pw_x_r = 20;
            32'b????_????_??10_0000_0000_0000_0000_0000:    Pw_x_r = 21;
            32'b????_????_?100_0000_0000_0000_0000_0000:    Pw_x_r = 22;
            32'b????_????_1000_0000_0000_0000_0000_0000:    Pw_x_r = 23;

            32'b????_???1_0000_0000_0000_0000_0000_0000:    Pw_x_r = 24;
            32'b????_??10_0000_0000_0000_0000_0000_0000:    Pw_x_r = 25;
            32'b????_?100_0000_0000_0000_0000_0000_0000:    Pw_x_r = 26;
            32'b????_1000_0000_0000_0000_0000_0000_0000:    Pw_x_r = 27;
            32'b???1_0000_0000_0000_0000_0000_0000_0000:    Pw_x_r = 28;
            32'b??10_0000_0000_0000_0000_0000_0000_0000:    Pw_x_r = 29;
            32'b?100_0000_0000_0000_0000_0000_0000_0000:    Pw_x_r = 30;
            32'b1000_0000_0000_0000_0000_0000_0000_0000:    Pw_x_r = 31;
            default:                                        Pw_x_r = 0;
        endcase

        casez (free_list_y)
            32'b????_????_????_????_????_????_????_???1:    Pw_y_r = 0;
            32'b????_????_????_????_????_????_????_??10:    Pw_y_r = 1;
            32'b????_????_????_????_????_????_????_?100:    Pw_y_r = 2;
            32'b????_????_????_????_????_????_????_1000:    Pw_y_r = 3;
            32'b????_????_????_????_????_????_???1_0000:    Pw_y_r = 4;
            32'b????_????_????_????_????_????_??10_0000:    Pw_y_r = 5;
            32'b????_????_????_????_????_????_?100_0000:    Pw_y_r = 6;
            32'b????_????_????_????_????_????_1000_0000:    Pw_y_r = 7;

            32'b????_????_????_????_????_???1_0000_0000:    Pw_y_r = 8;
            32'b????_????_????_????_????_??10_0000_0000:    Pw_y_r = 9;
            32'b????_????_????_????_????_?100_0000_0000:    Pw_y_r = 10;
            32'b????_????_????_????_????_1000_0000_0000:    Pw_y_r = 11;
            32'b????_????_????_????_???1_0000_0000_0000:    Pw_y_r = 12;
            32'b????_????_????_????_??10_0000_0000_0000:    Pw_y_r = 13;
            32'b????_????_????_????_?100_0000_0000_0000:    Pw_y_r = 14;
            32'b????_????_????_????_1000_0000_0000_0000:    Pw_y_r = 15;

            32'b????_????_????_???1_0000_0000_0000_0000:    Pw_y_r = 16;
            32'b????_????_????_??10_0000_0000_0000_0000:    Pw_y_r = 17;
            32'b????_????_????_?100_0000_0000_0000_0000:    Pw_y_r = 18;
            32'b????_????_????_1000_0000_0000_0000_0000:    Pw_y_r = 19;
            32'b????_????_???1_0000_0000_0000_0000_0000:    Pw_y_r = 20;
            32'b????_????_??10_0000_0000_0000_0000_0000:    Pw_y_r = 21;
            32'b????_????_?100_0000_0000_0000_0000_0000:    Pw_y_r = 22;
            32'b????_????_1000_0000_0000_0000_0000_0000:    Pw_y_r = 23;

            32'b????_???1_0000_0000_0000_0000_0000_0000:    Pw_y_r = 24;
            32'b????_??10_0000_0000_0000_0000_0000_0000:    Pw_y_r = 25;
            32'b????_?100_0000_0000_0000_0000_0000_0000:    Pw_y_r = 26;
            32'b????_1000_0000_0000_0000_0000_0000_0000:    Pw_y_r = 27;
            32'b???1_0000_0000_0000_0000_0000_0000_0000:    Pw_y_r = 28;
            32'b??10_0000_0000_0000_0000_0000_0000_0000:    Pw_y_r = 29;
            32'b?100_0000_0000_0000_0000_0000_0000_0000:    Pw_y_r = 30;
            32'b1000_0000_0000_0000_0000_0000_0000_0000:    Pw_y_r = 31;
            default:                                        Pw_y_r = 0;
        endcase

        casez (free_list_z)
            32'b????_????_????_????_????_????_????_???1:    Pw_z_r = 0;
            32'b????_????_????_????_????_????_????_??10:    Pw_z_r = 1;
            32'b????_????_????_????_????_????_????_?100:    Pw_z_r = 2;
            32'b????_????_????_????_????_????_????_1000:    Pw_z_r = 3;
            32'b????_????_????_????_????_????_???1_0000:    Pw_z_r = 4;
            32'b????_????_????_????_????_????_??10_0000:    Pw_z_r = 5;
            32'b????_????_????_????_????_????_?100_0000:    Pw_z_r = 6;
            32'b????_????_????_????_????_????_1000_0000:    Pw_z_r = 7;

            32'b????_????_????_????_????_???1_0000_0000:    Pw_z_r = 8;
            32'b????_????_????_????_????_??10_0000_0000:    Pw_z_r = 9;
            32'b????_????_????_????_????_?100_0000_0000:    Pw_z_r = 10;
            32'b????_????_????_????_????_1000_0000_0000:    Pw_z_r = 11;
            32'b????_????_????_????_???1_0000_0000_0000:    Pw_z_r = 12;
            32'b????_????_????_????_??10_0000_0000_0000:    Pw_z_r = 13;
            32'b????_????_????_????_?100_0000_0000_0000:    Pw_z_r = 14;
            32'b????_????_????_????_1000_0000_0000_0000:    Pw_z_r = 15;

            32'b????_????_????_???1_0000_0000_0000_0000:    Pw_z_r = 16;
            32'b????_????_????_??10_0000_0000_0000_0000:    Pw_z_r = 17;
            32'b????_????_????_?100_0000_0000_0000_0000:    Pw_z_r = 18;
            32'b????_????_????_1000_0000_0000_0000_0000:    Pw_z_r = 19;
            32'b????_????_???1_0000_0000_0000_0000_0000:    Pw_z_r = 20;
            32'b????_????_??10_0000_0000_0000_0000_0000:    Pw_z_r = 21;
            32'b????_????_?100_0000_0000_0000_0000_0000:    Pw_z_r = 22;
            32'b????_????_1000_0000_0000_0000_0000_0000:    Pw_z_r = 23;

            32'b????_???1_0000_0000_0000_0000_0000_0000:    Pw_z_r = 24;
            32'b????_??10_0000_0000_0000_0000_0000_0000:    Pw_z_r = 25;
            32'b????_?100_0000_0000_0000_0000_0000_0000:    Pw_z_r = 26;
            32'b????_1000_0000_0000_0000_0000_0000_0000:    Pw_z_r = 27;
            32'b???1_0000_0000_0000_0000_0000_0000_0000:    Pw_z_r = 28;
            32'b??10_0000_0000_0000_0000_0000_0000_0000:    Pw_z_r = 29;
            32'b?100_0000_0000_0000_0000_0000_0000_0000:    Pw_z_r = 30;
            32'b1000_0000_0000_0000_0000_0000_0000_0000:    Pw_z_r = 31;
            default:                                        Pw_z_r = 0;
        endcase
    end

    assign  full_PRF_x = (free_list == 32'd0)? 1 : 0;
    assign  full_PRF_y = (free_list_y == 32'd0)? 1 : 0;
    assign  full_PRF_z = (free_list_z == 32'd0)? 1 : 0;
    assign  full_PRF = (full_PRF_x || full_PRF_y || full_PRF_z)? 1 : 0;

endmodule