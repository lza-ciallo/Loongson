module PC (
    input               clk,
    input               rst,
    input               freeze_front,
    output  [7 : 0]     pc,
    output              valid_pc
);

endmodule