module DECODER (
    input   [9 : 0]     inst,
    output  [2 : 0]     Ra,
    output  [2 : 0]     Rb,
    output  [2 : 0]     Rw,
    input               valid_pc,
    output              valid_add,
    output              valid_mul
);

endmodule