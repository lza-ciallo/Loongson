// 最基本设定
