module PC (
    input clk,
    input rst,
    output [31:0] pc,
    input stall,
    // PC RENEW
    input jump,
    input [31:0] pc_jump,
    input predict,
    input [31:0] pc_predict,
    input rewind,
    input [31:0] pc_unsel
);




endmodule
