//
// IF 

`ifndef DEFINE
`define DEFINE
