module INST_MEM (
    input               rst,
    input   [7 : 0]     pc,
    output  [9 : 0]     inst_x,
    output  [9 : 0]     inst_y,
    output  [9 : 0]     inst_z
);

endmodule