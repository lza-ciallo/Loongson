`define     INT     5'b0000_0
`define     ADEF    5'b1000_0
`define     ADEM    5'b1000_1
`define     ALE     5'b1001_0
`define     SYS     5'b1011_0
`define     BRK     5'b1100_0
`define     INE     5'b1101_0
`define     IPE     5'b1110_0