// ALU
`define     ADD     32'b0000_0000_0001_0000_0???_????_????_????
`define     SUB     32'b0000_0000_0001_0001_0???_????_????_????
`define     SLT     32'b0000_0000_0001_0010_0???_????_????_????
`define     SLTU    32'b0000_0000_0001_0010_1???_????_????_????
`define     NOR     32'b0000_0000_0001_0100_0???_????_????_????
`define     AND     32'b0000_0000_0001_0100_1???_????_????_????
`define     OR      32'b0000_0000_0001_0101_0???_????_????_????
`define     XOR     32'b0000_0000_0001_0101_1???_????_????_????
`define     SLL     32'b0000_0000_0001_0111_0???_????_????_????
`define     SRL     32'b0000_0000_0001_0111_1???_????_????_????
`define     SRA     32'b0000_0000_0001_1000_0???_????_????_????

`define     SLLI    32'b0000_0000_0100_0000_1???_????_????_????
`define     SRLI    32'b0000_0000_0100_0100_1???_????_????_????
`define     SRAI    32'b0000_0000_0100_1000_1???_????_????_????

`define     SLTI    32'b0000_0010_00??_????_????_????_????_????
`define     SLTUI   32'b0000_0010_01??_????_????_????_????_????
`define     ADDI    32'b0000_0010_10??_????_????_????_????_????
`define     ANDI    32'b0000_0011_01??_????_????_????_????_????
`define     ORI     32'b0000_0011_10??_????_????_????_????_????
`define     XORI    32'b0000_0011_11??_????_????_????_????_????

// MDU
`define     MUL     32'b0000_0000_0001_1100_0???_????_????_????
`define     MULH    32'b0000_0000_0001_1100_1???_????_????_????
`define     MULHU   32'b0000_0000_0001_1101_0???_????_????_????
`define     DIV     32'b0000_0000_0010_0000_0???_????_????_????
`define     MOD     32'b0000_0000_0010_0000_1???_????_????_????
`define     DIVU    32'b0000_0000_0010_0001_0???_????_????_????
`define     MODU    32'b0000_0000_0010_0001_1???_????_????_????

// LSU
`define     LDB     32'b0010_1000_00??_????_????_????_????_????
`define     LDH     32'b0010_1000_01??_????_????_????_????_????
`define     LDW     32'b0010_1000_10??_????_????_????_????_????
`define     STB     32'b0010_1001_00??_????_????_????_????_????
`define     STH     32'b0010_1001_01??_????_????_????_????_????
`define     STW     32'b0010_1001_10??_????_????_????_????_????
`define     LDBU    32'b0010_1010_00??_????_????_????_????_????
`define     LDHU    32'b0010_1010_01??_????_????_????_????_????

// BRU
`define     BEQ     32'b0101_10??_????_????_????_????_????_????
`define     BNE     32'b0101_11??_????_????_????_????_????_????
`define     BLT     32'b0110_00??_????_????_????_????_????_????
`define     BGE     32'b0110_01??_????_????_????_????_????_????
`define     BLTU    32'b0110_10??_????_????_????_????_????_????
`define     BGEU    32'b0110_11??_????_????_????_????_????_????
`define     JIRL    32'b0100_11??_????_????_????_????_????_????

// DIR
`define     B       32'b0101_00??_????_????_????_????_????_????
`define     BL      32'b0101_01??_????_????_????_????_????_????
`define     LU12I   32'b0001_010?_????_????_????_????_????_????
`define     PCADD   32'b0001_110?_????_????_????_????_????_????

`define     CNTID   32'b0000_0000_0000_0000_0110_00??_???0_0000
`define     CNTVL   32'b0000_0000_0000_0000_0110_0000_000?_????
`define     CNTVH   32'b0000_0000_0000_0000_0110_0100_000?_????
`define     BREAK   32'b0000_0000_0010_1010_0???_????_????_????
`define     SYSCL   32'b0000_0000_0010_1011_0???_????_????_????

`define     CSR3    32'b0000_0100_????_????_????_????_????_????
`define     ERTN    32'b0000_0110_0100_1000_0011_1000_0000_0000
`define     IDLE    32'b0000_0110_0100_1000_1???_????_????_????

// 不打算实现
`define     CACOP   32'b0000_0110_00??_????_????_????_????_????
`define     TLBSH   32'b0000_0110_0100_1000_0010_1000_0000_0000
`define     TLBRD   32'b0000_0110_0100_1000_0010_1100_0000_0000
`define     TLBWR   32'b0000_0110_0100_1000_0011_0000_0000_0000
`define     TLBFL   32'b0000_0110_0100_1000_0011_0100_0000_0000
`define     INVTLB  32'b0000_0110_0100_1001_1???_????_????_????

`define     LL      32'b0010_0000_????_????_????_????_????_????
`define     SC      32'b0010_0001_????_????_????_????_????_????
`define     PRELD   32'b0010_1010_11??_????_????_????_????_????
`define     DBAR    32'b0011_1000_0111_0010_0???_????_????_????
`define     IBAR    32'b0011_1000_0111_0010_1???_????_????_????

`define     NOP     32'b0000_0000_0000_0000_0000_0000_0000_0000