module inst_mem (
    input               clk,
    input   [31 : 0]    pc,
    output  [31 : 0]    inst    [2 : 0]
);

    // 实例化一个 BRAM

endmodule